`default_nettype none

module uart_to_qspi (
    input wire clk,
    input wire resetn,
    // UART interface
    output wire ser_tx,
    input wire ser_rx,
    // QSPI interface
    input wire [3:0] qspi_io_in,    // 4-bit input from QSPI core
    output reg [3:0] qspi_io_out,   // 4-bit output to QSPI core
    output reg qspi_csb,            // Chip select (active low)
    output reg qspi_sck,            // Clock generated by bridge
    output reg [3:0] qspi_io_oe,    // Output enable FOR THE BRIDGE->CORE PATH
    // Management UART (unused in this setup)
    output wire mgmt_uart_rx,
    input wire mgmt_uart_tx,
    input wire mgmt_uart_enabled
);
    // Baud rate divider for 100MHz clock -> ~9600 baud
    localparam UART_DIVIDER = 16'd10417;
    localparam UART_HALF_DIVIDER = UART_DIVIDER / 2;

    // QSPI Clock Generation (e.g., 2MHz QSPI clock)
    localparam QSPI_CLK_CYCLES = 50;
    localparam QSPI_CLK_HALF_CYCLES = QSPI_CLK_CYCLES / 2;

    //============ UART Receiver Section (No changes needed here) ============//
    reg [3:0] recv_state;
    reg [15:0] recv_divcnt;
    // reg [7:0] recv_pattern; // Replaced by recv_shifter
    reg [7:0] recv_shifter; // Shift register for incoming bits
    reg [7:0] recv_buf_data; // Buffer for the completed byte
    reg recv_buf_valid;      // Flag indicating recv_buf_data is valid
    reg ser_rx_sync;
    reg ser_rx_sync_prev;

    always @(posedge clk) begin // Synchronizer
        if (!resetn) begin ser_rx_sync <= 1; ser_rx_sync_prev <= 1; end
        else begin ser_rx_sync_prev <= ser_rx_sync; ser_rx_sync <= ser_rx; end
    end
    wire ser_rx_falling_edge = ser_rx_sync_prev & !ser_rx_sync;

    always @(posedge clk) begin // UART RX FSM
        if (!resetn) begin /* resets */ recv_state <= 0; recv_divcnt <= 0; /* recv_pattern <= 0; */ recv_shifter <= 0; recv_buf_data <= 0; recv_buf_valid <= 0; end // Removed recv_pattern reset, added recv_shifter reset
        else begin
            // if (recv_buf_valid) recv_buf_valid <= 0; // REMOVED: Make valid flag sticky until consumed by QSPI FSM
            recv_divcnt <= recv_divcnt + 1;
            case (recv_state)
                0: if (ser_rx_falling_edge) begin recv_state <= 1; recv_divcnt <= 0; end else recv_divcnt <= 0; // Reset counter if staying idle
                1: if (recv_divcnt >= UART_HALF_DIVIDER) if (!ser_rx_sync) begin recv_state <= 2; recv_divcnt <= 0; recv_shifter <= 8'b0; end else recv_state <= 0; // Check start bit validity, reset shifter
                2: if (recv_divcnt >= UART_DIVIDER) begin recv_shifter <= {ser_rx_sync, recv_shifter[7:1]}; recv_divcnt <= 0; recv_state <= 3; end // Sample bit 0, shift into MSB, go to state 3
                // States 3-9 handled by default case
                10: if (recv_divcnt >= UART_DIVIDER) begin // Check stop bit
                        if (ser_rx_sync) begin // Stop bit should be high
                            recv_buf_data <= recv_shifter; recv_buf_valid <= 1; // Latch data from shifter, set valid flag
                            $display("UART_RX: Received Byte %h (from shifter %h) at %t", recv_shifter, recv_shifter, $time);
                        end else begin
                            $display("UART_RX: Framing Error! at %t", $time);
                            // Don't set recv_buf_valid on error
                        end
                        recv_state <= 0; recv_divcnt <= 0; // Go back to idle
                    end
                default: // Handles states 3 (bit 1) through 9 (bit 7)
                    if (recv_state >= 3 && recv_state <= 9) begin
                        if (recv_divcnt >= UART_DIVIDER) begin
                            recv_shifter <= {ser_rx_sync, recv_shifter[7:1]}; // Sample data bit, shift into MSB
                            recv_divcnt <= 0;
                            if (recv_state == 9) begin // If just sampled bit 7
                                recv_state <= 10; // Go check stop bit
                            end else begin
                                recv_state <= recv_state + 1; // Go sample next bit
                            end
                        end
                    end else begin
                        recv_state <= 0; // Should not happen, safety reset
                    end
            endcase
        end
    end

    assign ser_tx = mgmt_uart_enabled ? (mgmt_uart_tx & retn_pattern[0]) : retn_pattern[0];
    assign mgmt_uart_rx = ser_rx;

    //============ QSPI Communication Section ============//
    reg [3:0] send_state;
    localparam QSPI_IDLE      = 0;
    localparam QSPI_SEND_HI   = 1;
    localparam QSPI_WAIT_HI   = 2;
    localparam QSPI_SEND_LO   = 3;
    localparam QSPI_WAIT_LO   = 4;
    localparam QSPI_READ_WAIT_HI = 5;
    localparam QSPI_READ_HI   = 6;
    // Removed READ_WAIT_LO and READ_LO as they were combined into READ_HI logic

    reg [3:0] send_byte_cnt;
    reg [15:0] qspi_clk_divcnt;
    reg [7:0] send_buf_data;
    reg [7:0] recv_qspi_byte;

    // FIFO for buffering QSPI results before UART TX
    localparam FIFO_DEPTH_BITS = 2; // 2^2 = 4 entries
    localparam FIFO_DEPTH = 1 << FIFO_DEPTH_BITS;
    reg [7:0] fifo_mem [FIFO_DEPTH-1:0];
    reg [FIFO_DEPTH_BITS-1:0] fifo_wptr;
    reg [FIFO_DEPTH_BITS-1:0] fifo_rptr;
    reg [FIFO_DEPTH_BITS:0] fifo_count; // Can hold values 0 to FIFO_DEPTH
    wire fifo_empty = (fifo_count == 0);
    wire fifo_full = (fifo_count == FIFO_DEPTH);
    reg fifo_write_enable; // Pulse high for one cycle to write
    reg fifo_read_enable;  // Pulse high for one cycle to read
    wire [7:0] fifo_data_out = fifo_mem[fifo_rptr]; // Read directly from current rptr

    // QSPI return data communication (UART TX)
    reg [7:0] retn_buf_data; // Data currently being transmitted by UART
    // reg retn_req; // Replaced by FIFO empty check
    reg [3:0] retn_state;      // UART TX state machine
    reg [9:0] retn_pattern;
    reg [3:0] retn_bitcnt;
    reg [15:0] retn_divcnt;    // UART TX baud rate counter

    reg [3:0] result_counter;
    reg result_nibble_flag;

    always @(posedge clk) begin // QSPI FSM
        if (!resetn) begin
            qspi_clk_divcnt <= 0; send_state <= QSPI_IDLE; send_byte_cnt <= 0; send_buf_data <= 0;
            recv_qspi_byte <= 0; qspi_csb <= 1; qspi_sck <= 0; qspi_io_out <= 4'b0000; qspi_io_oe <= 4'b0000;
            // retn_req <= 0; // Removed retn_req
            result_counter <= 0; result_nibble_flag <= 0;

            // Reset FIFO
            fifo_wptr <= 0; fifo_rptr <= 0; fifo_count <= 0;
            fifo_write_enable <= 0; fifo_read_enable <= 0;

        end else begin
            // Default FIFO control signals (pulsed high when needed)
            fifo_write_enable <= 0;
            fifo_read_enable <= 0;

            qspi_clk_divcnt <= qspi_clk_divcnt + 1; // Advance QSPI clock divider

            // State transitions now based on QSPI clock timing derived from qspi_clk_divcnt
            case (send_state)
                QSPI_IDLE: begin
                    qspi_sck <= 0; qspi_clk_divcnt <= 0; qspi_io_oe <= 4'b0000;
                    if (recv_buf_valid) begin // Check if first byte is ready
                        recv_buf_valid <= 0; // Consume the byte
                        qspi_csb <= 0; send_state <= QSPI_SEND_HI; send_byte_cnt <= 0; send_buf_data <= recv_buf_data;
                        qspi_clk_divcnt <= 0; qspi_io_oe <= 4'b1111; qspi_io_out <= recv_buf_data[7:4]; qspi_sck <= 0;
                        $display("QSPI: Starting transaction, sending byte 0: %h at %t", recv_buf_data, $time);
                    end
                end

                QSPI_SEND_HI: begin // Wait half QSPI clock, raise clock
                    if (qspi_clk_divcnt >= QSPI_CLK_HALF_CYCLES) begin
                        qspi_sck <= 1; send_state <= QSPI_WAIT_HI; qspi_clk_divcnt <= 0;
                    end
                end

                QSPI_WAIT_HI: begin // Wait half QSPI clock, lower clock, prepare low nibble
                    if (qspi_clk_divcnt >= QSPI_CLK_HALF_CYCLES) begin
                        qspi_sck <= 0; qspi_io_out <= send_buf_data[3:0]; send_state <= QSPI_SEND_LO; qspi_clk_divcnt <= 0;
                    end
                end

                QSPI_SEND_LO: begin // Wait half QSPI clock, raise clock
                    if (qspi_clk_divcnt >= QSPI_CLK_HALF_CYCLES) begin
                        qspi_sck <= 1; send_state <= QSPI_WAIT_LO; qspi_clk_divcnt <= 0;
                    end
                end

                QSPI_WAIT_LO: begin // Wait half QSPI clock, lower clock, check if more bytes
                    if (qspi_clk_divcnt >= QSPI_CLK_HALF_CYCLES) begin
                        qspi_sck <= 0; qspi_clk_divcnt <= 0;
                        if (send_byte_cnt == 7) begin
                            $display("QSPI: Sent 8 bytes, moving to read results at %t", $time);
                            send_state <= QSPI_READ_WAIT_HI; qspi_io_oe <= 4'b0000;
                            result_counter <= 0; result_nibble_flag <= 0;
                        end else begin // Need to send more bytes (1-7)
                            if (recv_buf_valid) begin // Check if next UART byte is ready
                                recv_buf_valid <= 0; // Consume the byte
                                send_byte_cnt <= send_byte_cnt + 1; send_buf_data <= recv_buf_data;
                                qspi_io_out <= recv_buf_data[7:4]; send_state <= QSPI_SEND_HI;
                                $display("QSPI: Sending byte %d: %h at %t", send_byte_cnt + 1, recv_buf_data, $time);
                            end else begin
                                // Stay in QSPI_WAIT_LO, waiting for UART data
                                $display("QSPI: Waiting for sticky UART byte %d... at %t", send_byte_cnt + 1, $time);
                            end
                        end
                    end
                end

                QSPI_READ_WAIT_HI: begin // Keep clock low, wait half cycle
                    qspi_io_oe <= 4'b0000; qspi_sck <= 0;
                    if (qspi_clk_divcnt >= QSPI_CLK_HALF_CYCLES) begin
                         qspi_sck <= 1; send_state <= QSPI_READ_HI; qspi_clk_divcnt <= 0;
                    end
                end

                QSPI_READ_HI: begin // Clock is high, core puts data. Wait half cycle, read on falling edge.
                    if (qspi_clk_divcnt >= QSPI_CLK_HALF_CYCLES) begin
                        if (!result_nibble_flag) begin
                            recv_qspi_byte[7:4] <= qspi_io_in; result_nibble_flag <= 1;
                            $display("RESULT: Received high nibble %h for result %d at %t", qspi_io_in, result_counter, $time);
                        end else begin
                            recv_qspi_byte[3:0] <= qspi_io_in; result_nibble_flag <= 0;
                            $display("RESULT: Received low nibble %h, complete byte %h for result %d at %t", qspi_io_in, {recv_qspi_byte[7:4], qspi_io_in}, result_counter, $time);
                            // retn_buf_data <= {recv_qspi_byte[7:4], qspi_io_in}; // Store in FIFO instead
                            // retn_req <= 1; // Write to FIFO instead
                            if (!fifo_full) begin
                                fifo_write_enable <= 1; // Pulse high to write to FIFO
                                $display("FIFO: Writing byte %h (result %d) at %t", {recv_qspi_byte[7:4], qspi_io_in}, result_counter, $time);
                            end else begin
                                $display("FIFO: ERROR - FIFO Full! Cannot write result %d at %t", result_counter, $time);
                                // Handle error? For now, just drop data if full.
                            end

                            if (result_counter == 3) begin
                                $display("QSPI: Read all 4 results. Deasserting CS. FIFO count: %d. at %t", fifo_count + (fifo_write_enable && !fifo_full), $time); // Adjust count display for current write
                                send_state <= QSPI_IDLE; qspi_csb <= 1; qspi_sck <= 0;
                            end else begin
                                result_counter <= result_counter + 1; // Increment for next byte
                                // Need to go back to READ_WAIT_HI for the next byte
                                send_state <= QSPI_READ_WAIT_HI;
                            end
                        end // End of 'else' for low nibble read

                        // Common logic for both nibbles: Lower clock, reset divider
                        qspi_sck <= 0; // Lower the clock
                        qspi_clk_divcnt <= 0; // Reset divider for next half cycle

                        // State transition is now handled within the if/else based on result_counter
                        // If result_counter was 3, state is already set to QSPI_IDLE.
                        // If result_counter < 3, state is already set back to QSPI_READ_WAIT_HI.
                        // No need for the unconditional 'send_state <= QSPI_READ_WAIT_HI;' here anymore.
                    end
                end
                default: send_state <= QSPI_IDLE;
            endcase
        end
    end

    //============ FIFO Logic ============//
    always @(posedge clk) begin
        if (!resetn) begin
            // Reset handled in main FSM reset block
            // Initialize memory? Optional, depends on synthesis tool.
        end else begin
            if (fifo_write_enable && !fifo_full) begin
                fifo_mem[fifo_wptr] <= {recv_qspi_byte[7:4], qspi_io_in}; // Data comes from QSPI reader
                fifo_wptr <= fifo_wptr + 1;
                fifo_count <= fifo_count + 1;
            end
            if (fifo_read_enable && !fifo_empty) begin
                // data_out is assigned combinationally: fifo_data_out = fifo_mem[fifo_rptr];
                fifo_rptr <= fifo_rptr + 1;
                fifo_count <= fifo_count - 1;
            end
        end
    end

    //============ UART Return Data Section ============//
    always @(posedge clk) begin
        if (!resetn) begin
            retn_pattern <= 10'b1111111111; retn_bitcnt <= 0; retn_divcnt <= 0; retn_state <= 0;
            // FIFO reset handled in main FSM reset block
        end else begin
            case (retn_state)
                0: begin // IDLE_TX
                    retn_pattern[0] <= 1'b1; // Keep line high
                    if (!fifo_empty) begin // Start transmission if FIFO has data
                        fifo_read_enable <= 1; // Pulse high to read from FIFO
                        retn_buf_data <= fifo_data_out; // Latch data from FIFO output
                        $display("FIFO: Reading byte %h for UART TX at %t. FIFO count before read: %d", fifo_data_out, fifo_count, $time);
                        retn_pattern <= {1'b1, fifo_data_out, 1'b0}; // Load shifter: Stop(1), Data(8), Start(0)
                        retn_bitcnt <= 10;
                        retn_divcnt <= 0;
                        retn_state <= 1;
                        $display("UART_TX: Starting transmission of %h at %t", fifo_data_out, $time);
                    end else begin
                         retn_divcnt <= 0; // Stay idle, reset counter
                    end
                end
                1: begin // SENDING_BITS
                    retn_divcnt <= retn_divcnt + 1;
                    if (retn_divcnt >= UART_DIVIDER) begin
                        retn_divcnt <= 0;
                        retn_pattern <= {1'b1, retn_pattern[9:1]}; // Shift out LSB (pattern[0])
                        retn_bitcnt <= retn_bitcnt - 1;
                        if (retn_bitcnt == 0) begin
                            retn_state <= 0; // Transmission complete
                            $display("UART_TX: Transmission complete at %t", $time);
                        end
                    end
                end
                default: retn_state <= 0;
            endcase
        end
    end

endmodule
`default_nettype wire
